* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT RCA gnd B3 B0 C0 A3 A0 vdd A2 A1 B2 B1 S3 S0 C4 S2 S1
** N=95 EP=16 IP=0 FDC=168
M0 35 A3 15 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=12680 $Y=2200 $D=0
M1 36 A0 16 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=12680 $Y=12370 $D=0
M2 gnd B3 35 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=13370 $Y=2200 $D=0
M3 gnd B0 36 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=13370 $Y=12370 $D=0
M4 41 B3 13 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=14870 $Y=2200 $D=0
M5 42 B0 14 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=14870 $Y=12370 $D=0
M6 gnd 6 41 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=15560 $Y=2200 $D=0
M7 gnd C0 42 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=15560 $Y=12370 $D=0
M8 37 A3 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=15940 $Y=-6405 $D=0
M9 gnd 37 43 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=15940 $Y=-4395 $D=0
M10 43 B3 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15940 $Y=-3705 $D=0
M11 4 39 43 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15940 $Y=-3015 $D=0
M12 43 A3 4 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=15940 $Y=-2325 $D=0
M13 gnd B3 39 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=15940 $Y=-305 $D=0
M14 40 B0 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=15940 $Y=15195 $D=0
M15 5 A0 44 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=15940 $Y=17215 $D=0
M16 44 40 5 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15940 $Y=17905 $D=0
M17 gnd B0 44 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15940 $Y=18595 $D=0
M18 44 38 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=15940 $Y=19285 $D=0
M19 gnd A0 38 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=15940 $Y=21295 $D=0
M20 45 6 8 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17060 $Y=2200 $D=0
M21 46 C0 9 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17060 $Y=12370 $D=0
M22 gnd A3 45 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=17750 $Y=2200 $D=0
M23 gnd A0 46 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=17750 $Y=12370 $D=0
M24 55 4 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=20060 $Y=-6405 $D=0
M25 gnd 55 47 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=20060 $Y=-4395 $D=0
M26 47 6 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20060 $Y=-3705 $D=0
M27 S3 51 47 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20060 $Y=-3015 $D=0
M28 47 4 S3 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=20060 $Y=-2325 $D=0
M29 gnd 6 51 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=20060 $Y=-305 $D=0
M30 54 C0 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=20060 $Y=15195 $D=0
M31 S0 5 48 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=20060 $Y=17215 $D=0
M32 48 54 S0 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20060 $Y=17905 $D=0
M33 gnd C0 48 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20060 $Y=18595 $D=0
M34 48 56 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=20060 $Y=19285 $D=0
M35 gnd 5 56 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=20060 $Y=21295 $D=0
M36 52 8 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=22395 $Y=2660 $D=0
M37 53 9 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=22395 $Y=11910 $D=0
M38 61 13 52 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23085 $Y=2660 $D=0
M39 62 14 53 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23085 $Y=11910 $D=0
M40 C4 15 61 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=23775 $Y=2660 $D=0
M41 18 16 62 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=23775 $Y=11910 $D=0
M42 68 29 6 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=27905 $Y=2660 $D=0
M43 69 30 17 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=27905 $Y=11910 $D=0
M44 70 25 68 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=28595 $Y=2660 $D=0
M45 71 26 69 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=28595 $Y=11910 $D=0
M46 gnd 19 70 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=29285 $Y=2660 $D=0
M47 gnd 20 71 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=29285 $Y=11910 $D=0
M48 72 21 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=31300 $Y=-6405 $D=0
M49 gnd 72 78 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=31300 $Y=-4395 $D=0
M50 78 17 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31300 $Y=-3705 $D=0
M51 S2 74 78 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31300 $Y=-3015 $D=0
M52 78 21 S2 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=31300 $Y=-2325 $D=0
M53 gnd 17 74 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=31300 $Y=-305 $D=0
M54 75 18 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=31300 $Y=15195 $D=0
M55 S1 22 79 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=31300 $Y=17215 $D=0
M56 79 75 S1 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31300 $Y=17905 $D=0
M57 gnd 18 79 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31300 $Y=18595 $D=0
M58 79 73 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=31300 $Y=19285 $D=0
M59 gnd 22 73 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=31300 $Y=21295 $D=0
M60 80 A2 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=33930 $Y=2200 $D=0
M61 81 A1 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=33930 $Y=12370 $D=0
M62 19 17 80 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=34620 $Y=2200 $D=0
M63 20 18 81 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=34620 $Y=12370 $D=0
M64 88 A2 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=35420 $Y=-6405 $D=0
M65 gnd 88 82 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=35420 $Y=-4395 $D=0
M66 82 B2 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=35420 $Y=-3705 $D=0
M67 21 86 82 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=35420 $Y=-3015 $D=0
M68 82 A2 21 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=35420 $Y=-2325 $D=0
M69 gnd B2 86 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=35420 $Y=-305 $D=0
M70 87 B1 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=35420 $Y=15195 $D=0
M71 22 A1 83 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=35420 $Y=17215 $D=0
M72 83 87 22 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=35420 $Y=17905 $D=0
M73 gnd B1 83 gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=35420 $Y=18595 $D=0
M74 83 89 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=35420 $Y=19285 $D=0
M75 gnd A1 89 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=35420 $Y=21295 $D=0
M76 84 17 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=36120 $Y=2200 $D=0
M77 85 18 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=36120 $Y=12370 $D=0
M78 25 B2 84 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=36810 $Y=2200 $D=0
M79 26 B1 85 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=36810 $Y=12370 $D=0
M80 90 B2 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=38310 $Y=2200 $D=0
M81 91 B1 gnd gnd N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=38310 $Y=12370 $D=0
M82 29 A2 90 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=39000 $Y=2200 $D=0
M83 30 A1 91 gnd N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=39000 $Y=12370 $D=0
M84 37 A3 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=12355 $Y=-6405 $D=1
M85 31 37 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=12355 $Y=-4395 $D=1
M86 4 B3 31 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=12355 $Y=-3705 $D=1
M87 32 39 4 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=12355 $Y=-3015 $D=1
M88 vdd A3 32 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=12355 $Y=-2325 $D=1
M89 vdd B3 39 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=12355 $Y=-305 $D=1
M90 40 B0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=12355 $Y=15195 $D=1
M91 33 A0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=12355 $Y=17215 $D=1
M92 5 40 33 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=12355 $Y=17905 $D=1
M93 34 B0 5 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=12355 $Y=18595 $D=1
M94 vdd 38 34 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=12355 $Y=19285 $D=1
M95 vdd A0 38 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=12355 $Y=21295 $D=1
M96 15 A3 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=12680 $Y=4285 $D=1
M97 16 A0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=12680 $Y=9785 $D=1
M98 vdd B3 15 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=13370 $Y=4285 $D=1
M99 vdd B0 16 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=13370 $Y=9785 $D=1
M100 13 B3 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=14870 $Y=4285 $D=1
M101 14 B0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=14870 $Y=9785 $D=1
M102 vdd 6 13 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=15560 $Y=4285 $D=1
M103 vdd C0 14 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=15560 $Y=9785 $D=1
M104 8 6 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17060 $Y=4285 $D=1
M105 9 C0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17060 $Y=9785 $D=1
M106 vdd A3 8 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=17750 $Y=4285 $D=1
M107 vdd A0 9 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=17750 $Y=9785 $D=1
M108 C4 8 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=22395 $Y=5050 $D=1
M109 18 9 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=22395 $Y=9020 $D=1
M110 vdd 13 C4 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23085 $Y=5050 $D=1
M111 vdd 14 18 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23085 $Y=9020 $D=1
M112 55 4 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=23145 $Y=-6405 $D=1
M113 57 55 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=23145 $Y=-4395 $D=1
M114 S3 6 57 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23145 $Y=-3705 $D=1
M115 58 51 S3 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23145 $Y=-3015 $D=1
M116 vdd 4 58 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=23145 $Y=-2325 $D=1
M117 vdd 6 51 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=23145 $Y=-305 $D=1
M118 54 C0 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=23145 $Y=15195 $D=1
M119 59 5 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=23145 $Y=17215 $D=1
M120 S0 54 59 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23145 $Y=17905 $D=1
M121 60 C0 S0 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=23145 $Y=18595 $D=1
M122 vdd 56 60 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=23145 $Y=19285 $D=1
M123 vdd 5 56 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=23145 $Y=21295 $D=1
M124 C4 15 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=23775 $Y=5050 $D=1
M125 18 16 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=23775 $Y=9020 $D=1
M126 72 21 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=27715 $Y=-6405 $D=1
M127 64 72 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=27715 $Y=-4395 $D=1
M128 S2 17 64 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=27715 $Y=-3705 $D=1
M129 65 74 S2 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=27715 $Y=-3015 $D=1
M130 vdd 21 65 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=27715 $Y=-2325 $D=1
M131 vdd 17 74 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=27715 $Y=-305 $D=1
M132 75 18 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=27715 $Y=15195 $D=1
M133 66 22 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=27715 $Y=17215 $D=1
M134 S1 75 66 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=27715 $Y=17905 $D=1
M135 67 18 S1 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=27715 $Y=18595 $D=1
M136 vdd 73 67 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=27715 $Y=19285 $D=1
M137 vdd 22 73 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=27715 $Y=21295 $D=1
M138 vdd 29 6 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=27905 $Y=5050 $D=1
M139 vdd 30 17 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=27905 $Y=9020 $D=1
M140 6 25 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=28595 $Y=5050 $D=1
M141 17 26 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=28595 $Y=9020 $D=1
M142 vdd 19 6 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=29285 $Y=5050 $D=1
M143 vdd 20 17 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=29285 $Y=9020 $D=1
M144 19 A2 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=33930 $Y=4285 $D=1
M145 20 A1 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=33930 $Y=9785 $D=1
M146 vdd 17 19 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=34620 $Y=4285 $D=1
M147 vdd 18 20 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=34620 $Y=9785 $D=1
M148 25 17 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=36120 $Y=4285 $D=1
M149 26 18 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=36120 $Y=9785 $D=1
M150 vdd B2 25 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=36810 $Y=4285 $D=1
M151 vdd B1 26 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=36810 $Y=9785 $D=1
M152 29 B2 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=38310 $Y=4285 $D=1
M153 30 B1 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=38310 $Y=9785 $D=1
M154 88 A2 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=38505 $Y=-6405 $D=1
M155 92 88 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=38505 $Y=-4395 $D=1
M156 21 B2 92 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=38505 $Y=-3705 $D=1
M157 93 86 21 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=38505 $Y=-3015 $D=1
M158 vdd A2 93 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=38505 $Y=-2325 $D=1
M159 vdd B2 86 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=38505 $Y=-305 $D=1
M160 87 B1 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=38505 $Y=15195 $D=1
M161 94 A1 vdd vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=38505 $Y=17215 $D=1
M162 22 87 94 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=38505 $Y=17905 $D=1
M163 95 B1 22 vdd P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=2.55e-13 PD=5.1e-07 PS=5.1e-07 $X=38505 $Y=18595 $D=1
M164 vdd 89 95 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=38505 $Y=19285 $D=1
M165 vdd A1 89 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=38505 $Y=21295 $D=1
M166 vdd A2 29 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=39000 $Y=4285 $D=1
M167 vdd A1 30 vdd P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07 $X=39000 $Y=9785 $D=1
.ENDS
***************************************
