**DFF**
.subckt DFF D CLK RESET Q QX VDD GND

**I1 I1vi1 I1vi2 I1vo VDD GND**
MpI1A	I1vo	I1vi1	VDD	VDD	p_18	W=1u	L=0.18u
MpI1B	I1vo	I1vi2	VDD	VDD	p_18	W=1u	L=0.18u
MnI1A2	I1vo	I1vi1	as1	GND	n_18	W=0.5u	L=0.18u
MnI1B2	as1	    I1vi2	GND	GND	n_18	W=0.5u	L=0.18u

**I2 I1vo CLK RESET I1vi2 VDD GND**
MpAI2  I1vi2 I1vo VDD  VDD p_18	W=1u	L=0.18u
MpBI2  I1vi2 CLK VDD  VDD p_18	W=1u	L=0.18u
MpCI2  I1vi2 RESET VDD  VDD p_18	W=1u	L=0.18u
MnAI22 I1vi2 I1vo as2  GND n_18	W=0.5u	L=0.18u
MnBI22 as2  CLK as22 GND n_18	W=0.5u	L=0.18u
MnCI22 as22 RESET GND  GND n_18	W=0.5u	L=0.18u

**I3 I1vi2 CLK I1vi1 I3vo VDD GND**
MpAI3  I3vo I1vi2 VDD  VDD p_18	W=1u	L=0.18u
MpBI3  I3vo CLK VDD  VDD p_18	W=1u	L=0.18u
MpCI3  I3vo I1vi1 VDD  VDD p_18	W=1u	L=0.18u
MnAI33 I3vo I1vi2 as3  GND n_18	W=0.5u	L=0.18u
MnBI33 as3  CLK as33 GND n_18	W=0.5u	L=0.18u
MnCI33 as33 I1vi1 GND  GND n_18	W=0.5u	L=0.18u

**I4 I3vo D RESET I1vi1 VDD GND**
MpAI4  I1vi1 I3vo VDD  VDD p_18	W=1u	L=0.18u
MpBI4  I1vi1 D VDD  VDD p_18	W=1u	L=0.18u
MpCI4  I1vi1 RESET VDD  VDD p_18	W=1u	L=0.18u
MnAI44 I1vi1 I3vo as4  GND n_18	W=0.5u	L=0.18u
MnBI44 as4  D as44 GND n_18	W=0.5u	L=0.18u
MnCI44 as44 RESET GND  GND n_18	W=0.5u	L=0.18u

**I5 I1vi2 QX Q VDD GND**
MpI5A	Q	I1vi2	VDD	VDD	p_18	W=1u	L=0.18u
MpI5B	Q	QX	VDD	VDD	p_18	W=1u	L=0.18u
MnI5A2	Q	I1vi2	as5	GND	n_18	W=0.5u	L=0.18u
MnI5B2	as5	    QX	GND	GND	n_18	W=0.5u	L=0.18u

**I6 Q I3vo RESET QX VDD GND**
MpAI6  QX Q VDD  VDD p_18	W=1u	L=0.18u
MpBI6  QX I3vo VDD  VDD p_18	W=1u	L=0.18u
MpCI6  QX RESET VDD  VDD p_18	W=1u	L=0.18u
MnAI66 QX Q as6  GND n_18	W=0.5u	L=0.18u
MnBI66 as6  I3vo as66 GND n_18	W=0.5u	L=0.18u
MnCI66 as66 RESET GND  GND n_18	W=0.5u	L=0.18u

.ends