***Lab12_RCA***
.include "fa.spi"

.subckt R_adder A0 B0 C0 A1 B1 A2 B2 A3 B3 C4 S0 S1 S2 S3 vdd gnd

	*fulladder 	A B C S COUT VDD GND
	Xfa1 A0 B0 C0 S0 C1 vdd gnd fulladder
	Xfa2 A1 B1 C1 S1 C2 vdd gnd fulladder
	Xfa3 A2 B2 C2 S2 C3 vdd gnd fulladder
	Xfa4 A3 B3 C3 S3 C4 vdd gnd fulladder

.ends